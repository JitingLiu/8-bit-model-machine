LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY model_machine IS
PORT(
	CLK_50M,CLR,rst: IN STD_LOGIC;
	clk_out: OUT STD_LOGIC;
	r_out,d_out: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	LD1,ADD1,SUB1,A_AND1,A_SRL1,HALT1:OUT STD_LOGIC;
	OUTPUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END model_machine;

ARCHITECTURE DATAFLOW OF model_machine IS
SIGNAL CLK,T0,T1,T2,T3,T4,T5,T6,T7: STD_LOGIC := '0';
SIGNAL LD,ADD,SUB,A_AND,A_SRL,HALT: STD_LOGIC := '0';
SIGNAL IPC,IMAR,IDR,EDR,IA,EA,ALU_ADD,ALU_SUB,ALU_AND,ALU_SRL,IIR: STD_LOGIC := '0'; --微指令输出
SIGNAL ACC_OUT,DR_OUT,ALU_OUT,RAM_OUT: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL PC_OUT,ADDR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
COMPONENT RAM IS 
PORT( 
	WR,CS:IN STD_LOGIC; --WR片选信号, CS读写控制端
	DIN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入的内存内容
	DOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --输出的是选中地址中相应的内容
	ADDR:IN STD_LOGIC_VECTOR(3 DOWNTO 0) ); --输入信号为地址信息
END COMPONENT; 

COMPONENT PC IS --程序计数器
PORT( 
	IPC,CLK,CLR:IN STD_LOGIC; 
	PCOUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0)  ); 
END COMPONENT;

COMPONENT MAR IS --保存当前 CPU 所访问的主存储器单元的地址
PORT( 
	ADDR_IN:IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
	IMAR:IN STD_LOGIC; 
	CLK:IN STD_LOGIC; 
	ADDR_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0) );
END COMPONENT;

COMPONENT IR IS --指令寄存器
PORT( 
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入
	IIR:IN STD_LOGIC; --使能。低有效
	CLK:IN STD_LOGIC; 
	LD,ADD,SUB,A_AND,A_SRL,HALT: OUT STD_LOGIC ); 
END COMPONENT;

COMPONENT DR IS --数据寄存器
PORT( 
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
	IDR:IN STD_LOGIC; 
	EDR:IN STD_LOGIC; 
	CLK:IN STD_LOGIC; 
	DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0) ); 
END COMPONENT;

COMPONENT COUNTER IS --节拍发生器
PORT( 
	CLK,CLR:IN STD_LOGIC; 
	T0,T1,T2,T3,T4,T5,T6,T7:OUT STD_LOGIC ); 
END COMPONENT;

COMPONENT CTRL IS --控制器
PORT( 
	LD,ADD,SUB,A_AND,A_SRL,HALT:IN STD_LOGIC; --操作指令信号
	CLK:IN STD_LOGIC; 
	T0,T1,T2,T3,T4,T5,T6,T7:IN STD_LOGIC; --节拍脉冲
	IPC,IMAR,IDR,EDR,IA,EA,ALU_ADD,ALU_SUB,ALU_AND,ALU_SRL,IIR:OUT STD_LOGIC ); --输出为十一个控制信号
END COMPONENT;

COMPONENT CLK_SOURCE IS
PORT(
	  CLK_50M:IN STD_LOGIC; 
	  CLK:OUT STD_LOGIC); --时钟周期为1s
END COMPONENT;

COMPONENT ALU IS
PORT(
 	rst:in std_logic;
  	acc:in std_logic_vector(7 downto 0);--累加器 	
	dr:in std_logic_vector(7 downto 0);--数据寄存器 		
	alu_add:in std_logic; --add加 	
	alu_sub:in std_logic; --sub减 	
	alu_and:in std_logic; --and与 	
	alu_srl:in std_logic; --srl左移 	
	alu_out:out std_logic_vector(7 downto 0)); --alu计算结果
END COMPONENT;

COMPONENT ACC IS
PORT( 
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入
	IA:IN STD_LOGIC; --输入控制信号
	EA:IN STD_LOGIC; --输出控制信号
	CLK:IN STD_LOGIC; 
	DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0) ); --输出
END COMPONENT;
BEGIN

M0: CLK_SOURCE PORT MAP (CLK_50M, CLK); --时钟例化
M1: COUNTER PORT MAP (CLK, CLR, T0, T1, T2, T3, T4, T5, T6, T7); --节拍例化
M2: CTRL PORT MAP (LD,ADD,SUB,A_AND,A_SRL,HALT,CLK,T0,T1,T2,T3,T4,T5,T6,T7, --控制器例化
						IPC,IMAR,IDR,EDR,IA,EA,ALU_ADD,ALU_SUB,ALU_AND,ALU_SRL,IIR); 
M3: ALU PORT MAP(rst,ACC_OUT,DR_OUT,ALU_ADD,ALU_SUB,ALU_AND,ALU_SRL,ALU_OUT); --算数逻辑单元
M4: ACC PORT MAP(DR_OUT, IA, EA, CLK, ACC_OUT); --累加器
M5: DR  PORT MAP(RAM_OUT, IDR, EDR, CLK, DR_OUT); --数据寄存器
M6: PC  PORT MAP(IPC,CLK,CLR,PC_OUT);
M7: MAR PORT MAP(PC_OUT,IMAR,CLK,ADDR_OUT); 
M8: IR  PORT MAP(DR_OUT,IIR,CLK,LD,ADD,SUB,A_AND,A_SRL,HALT); --指令寄存器
M9: RAM PORT MAP('1','0',"00000000",RAM_OUT,ADDR_OUT); --存储器
OUTPUT <= ALU_OUT;
r_out <= ACC_OUT;
d_out <= DR_OUT;
clk_out <= clk;
LD1<=LD; ADD1<=ADD; SUB1<=SUB; A_AND1<=A_AND; A_SRL1<=A_SRL; HALT1<=HALT;

END DATAFLOW;