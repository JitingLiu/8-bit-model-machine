LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
ENTITY MAR IS --保存当前 CPU 所访问的主存储器单元的地址
PORT( 
	ADDR_IN:IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
	IMAR:IN STD_LOGIC; 
	CLK:IN STD_LOGIC; 
	ADDR_OUT:OUT STD_LOGIC_VECTOR(3 DOWNTO 0) );
END MAR; 
 
ARCHITECTURE A OF MAR IS 
BEGIN 
	PROCESS(CLK,IMAR,ADDR_IN) 
	BEGIN 
	IF(CLK'EVENT AND CLK='1') THEN 
		IF(IMAR='0') THEN 
			ADDR_OUT<=ADDR_IN; 
		END IF; 
	END IF; 
	END PROCESS; 
END A;