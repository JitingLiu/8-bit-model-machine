LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
ENTITY IR IS --指令寄存器
PORT( 
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入
	IIR:IN STD_LOGIC; --使能。低有效
	CLK:IN STD_LOGIC; 
	LD,ADD,SUB,A_AND,A_SRL,HALT: OUT STD_LOGIC ); 
END IR; 

ARCHITECTURE DATAFLOW OF IR IS 
SIGNAL REGQ: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN 
	PROCESS(CLK,IIR) 
	BEGIN 
	IF(CLK'EVENT AND CLK='1') THEN 
		IF(IIR='0') THEN 
			REGQ<=DATA_IN; 
		END IF; 
	END IF; 
	END PROCESS; 
 
	PROCESS(CLK,REGQ) 
	BEGIN 
	CASE REGQ IS 
		WHEN "00111110" => LD<='1';ADD<='0';SUB<='0';A_AND<='0';A_SRL<='0';HALT<='0'; 
		WHEN "11000110" => LD<='0';ADD<='1';SUB<='0';A_AND<='0';A_SRL<='0';HALT<='0'; 
		WHEN "00110011" => LD<='0';ADD<='0';SUB<='1';A_AND<='0';A_SRL<='0';HALT<='0'; 
		WHEN "01110001" => LD<='0';ADD<='0';SUB<='0';A_AND<='1';A_SRL<='0';HALT<='0'; 
		WHEN "10110110" => LD<='0';ADD<='0';SUB<='0';A_AND<='0';A_SRL<='1';HALT<='0'; 
		WHEN "01110110" => LD<='0';ADD<='0';SUB<='0';A_AND<='0';A_SRL<='0';HALT<='1'; 
		WHEN OTHERS =>NULL; 
	END CASE; 
	END PROCESS; 
END DATAFLOW;