LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY CTRL IS 
	PORT( 
	LD,ADD,SUB,A_AND,A_SRL,HALT:IN STD_LOGIC; --操作指令信号
	CLK:IN STD_LOGIC; 
	T0,T1,T2,T3,T4,T5,T6,T7:IN STD_LOGIC; --节拍脉冲
	IPC,IMAR,IDR,EDR,IA,EA,ALU_ADD,ALU_SUB,ALU_AND,ALU_SRL,IIR:OUT STD_LOGIC ); --输出为十一个控制信号
END ENTITY; 

ARCHITECTURE A OF CTRL IS 
BEGIN 
	PROCESS(CLK,LD,ADD,SUB,A_AND,A_SRL,HALT,T0,T1,T2,T3,T4,T5,T6,T7) 
	BEGIN 
	IF(HALT='1')THEN 
		IPC<='0'; 	
	ELSE 
		IMAR<= NOT(T0 OR (T3 AND LD) OR (T3 AND ADD) OR (T3 AND SUB) OR (T3 AND A_AND) OR (T3 AND A_SRL)); 
		IIR <= NOT T2; 
		IA  <= NOT((T6 AND LD) OR (T6 AND ADD) OR (T6 AND SUB) OR (T6 AND A_AND) OR (T6 AND A_SRL)); 
		IDR <= T1 OR (T4 AND LD) OR (T4 AND ADD) OR (T4 AND SUB) OR (T4 AND A_AND) OR (T4 AND A_SRL); 
		IPC <= T2 OR (T5 AND LD) OR (T5 AND ADD) OR (T5 AND SUB) OR (T5 AND A_AND); 
		ALU_ADD <= NOT(T5 AND ADD); --加法
		ALU_SUB <= NOT(T5 AND SUB); --减法
		ALU_AND <= NOT(T5 AND A_AND); --与运算
		ALU_SRL <= NOT(T5 AND A_SRL); --左移
		EA <= '0';--(T7 AND ADD) OR (T7 AND SUB) OR (T7 AND A_AND) OR (T7 AND A_SRL); 
		EDR<= '0'; 
	END IF; 
	END PROCESS; 
END A;